.include TSMC_180nm.txt
.include subckt.txt

.param SUPPLY=1.8
.param LAMBDA = 0.09u
.param len = 2*LAMBDA
.param W_P = 20*LAMBDA
.param W_N = 10*LAMBDA

.global gnd vdd 
vdd vdd gnd 'SUPPLY'

* Input Pulses
VA A gnd pulse (0 SUPPLY 10ns .1ns .1ns 10ns 20ns)
VB B gnd pulse (0 SUPPLY 20ns .1ns .1ns 20ns 40ns)
* VC C gnd pulse (0 SUPPLY 40ns .1ns .1ns 40ns 80ns)
* VC D gnd pulse (0 SUPPLY 80ns .1ns .1ns 80ns 160ns)
VE en gnd pulse (0 SUPPLY 5ns .1ns .1ns 20ns 40ns)

* D-Latch Implementation

.subckt d_latch q d en vdd gnd 
Xinv d_inv d vdd gnd inv
Xnand1 out_n1 d en vdd gnd nand2
Xnand2 out_n2 d_inv en vdd gnd nand2
Xnand3 q out_n1 q1 vdd gnd nand2
Xnand4 q1 out_n2 q vdd gnd nand2
* Xbuff q_final q vdd gnd buffer
.ends d_latch

* Instantiate D-Latch
Xdlat q A en vdd gnd d_latch

* Simulation Setup
.tran 0.01ns 80ns
.control
    set hcopypscolor = 1
    set color0 = black
    set color1 = white
    run
    set curplottitle= d_latch
    plot v(A) v(en) v(q)+2
.endc
.end